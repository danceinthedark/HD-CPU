module HDCPU()
endmodule 